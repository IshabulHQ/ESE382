-------------------------------------------------------------------------------
--
-- Title       : gray_bin
-- Design      : gray_bin_csop
-- Author      : Ishabul Haque
-- Company     : stony brook
--
-------------------------------------------------------------------------------
--
-- File        : \\Mac\Home\Desktop\ESE382\Lab3\gray_to_binary\gray_bin_csop\src\gray_bin.vhd
-- Generated   : Tue Feb 18 23:47:28 2020
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {gray_bin} architecture {gray_bin}}

library IEEE;
use IEEE.std_logic_1164.all;

entity gray_bin is
	 port(
		 g3 : in STD_LOGIC;
		 g2 : in STD_LOGIC;
		 g1 : in STD_LOGIC;
		 g0 : in STD_LOGIC;
		 b3 : out STD_LOGIC;
		 b2 : out STD_LOGIC;
		 b1 : out STD_LOGIC;
		 b0 : out STD_LOGIC
	     );
end gray_bin;

--}} End of automatically maintained section

architecture gray_bin of gray_bin is
begin

	 -- enter your statements here --

end gray_bin;
